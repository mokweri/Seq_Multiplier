library verilog;
use verilog.vl_types.all;
entity Seq_Multiplier_tb is
end Seq_Multiplier_tb;
